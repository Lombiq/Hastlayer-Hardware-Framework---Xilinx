library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library Hast;
use Hast.SimpleMemory.all;

entity Hast_IP is 
    port(
        \DataIn\: In std_logic_vector(31 downto 0);
        \DataOut\: Out std_logic_vector(31 downto 0);
        \CellIndex\: Out integer;
        \ReadEnable\: Out boolean;
        \WriteEnable\: Out boolean;
        \ReadsDone\: In boolean;
        \WritesDone\: In boolean;
        \MemberId\: In integer;
        \Reset\: In std_logic;
        \Started\: In boolean;
        \Finished\: Out boolean;
        \Clock\: In std_logic
    );
    -- Hast_IP ID: -1989276552
    -- Date and time: 2016.07.23. 10:43:49 UTC
    -- Generated by Hastlayer - hastlayer.com
end Hast_IP;

architecture Imp of Hast_IP is 
    -- This IP was generated by Hastlayer from .NET code to mimic the original logic. Note the following:
    -- * For each member (methods, functions) in .NET a state machine was generated. Each state machine's name corresponds to 
    --   the original member's name.
    -- * Inputs and outputs are passed between state machines as shared objects.
    -- * There are operations that take multiple clock cycles like interacting with the memory and long-running arithmetic operations 
    --   (modulo, division, multiplication). These are awaited in subsequent states but be aware that some states can take more 
    --   than one clock cycle to produce their output.
    -- * The ExternalInvocationProxy process dispatches invocations that were started from the outside to the state machines.
    -- * The InternalInvocationProxy processes dispatch invocations between state machines.

    -- Array declarations start
    type boolean_Array is array (integer range <>) of boolean;
    -- Array declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).0 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).0 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).1 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).1 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).2 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).2 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).3 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).3 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).4 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).4 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).5 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).5 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).6 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).6 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).7 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).7 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).8 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).8 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).9 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).9 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).10 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).10 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).11 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).11 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).12 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).12 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).13 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).13 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).14 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).14 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).15 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).15 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).16 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).16 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).17 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).17 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).18 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).18 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).19 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).19 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).20 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).20 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).21 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).21 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).22 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).22 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).23 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).23 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).24 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).24 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).25 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).25 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).26 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).26 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).27 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).27 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).28 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).28 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).29 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).29 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).30 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).30 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).31 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).31 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).32 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).32 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).33 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).33 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).34 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.return\: boolean;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.numberObject.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).34 declarations end


    -- System.Void Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumber(Hast.Transformer.SimpleMemory.SimpleMemory).0 declarations start
    -- State machine states:
    type \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._States\ is (
        \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_0\, 
        \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_1\, 
        \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_2\, 
        \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_3\, 
        \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_4\, 
        \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_5\);
    -- Signals:
    Signal \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Finished\: boolean := false;
    Signal \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.CellIndex\: signed(31 downto 0);
    Signal \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.DataOut\: std_logic_vector(31 downto 0);
    Signal \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.ReadEnable\: boolean := false;
    Signal \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.WriteEnable\: boolean := false;
    Signal \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32).number.parameter.0\: unsigned(31 downto 0);
    Signal \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Started.0\: boolean := false;
    Signal \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Started\: boolean := false;
    Signal \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Finished.0\: boolean := false;
    Signal \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32).return.0\: boolean;
    -- System.Void Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumber(Hast.Transformer.SimpleMemory.SimpleMemory).0 declarations end


    -- System.Threading.Tasks.Task Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberAsync(Hast.Transformer.SimpleMemory.SimpleMemory).0 declarations start
    -- State machine states:
    type \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._States\ is (
        \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State_0\, 
        \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State_1\, 
        \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State_2\, 
        \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State_3\);
    -- Signals:
    Signal \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._Finished\: boolean := false;
    Signal \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.PrimeCalculator::IsPrimeNumber(SimpleMemory)._Started.0\: boolean := false;
    Signal \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._Started\: boolean := false;
    Signal \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.PrimeCalculator::IsPrimeNumber(SimpleMemory)._Finished.0\: boolean := false;
    -- System.Threading.Tasks.Task Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberAsync(Hast.Transformer.SimpleMemory.SimpleMemory).0 declarations end


    -- System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 declarations start
    -- State machine states:
    type \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._States\ is (
        \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_0\, 
        \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_1\, 
        \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_2\, 
        \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_3\, 
        \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_4\, 
        \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_5\, 
        \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_6\, 
        \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_7\, 
        \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_8\);
    -- Signals:
    Signal \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._Finished\: boolean := false;
    Signal \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.CellIndex\: signed(31 downto 0);
    Signal \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.DataOut\: std_logic_vector(31 downto 0);
    Signal \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\: boolean := false;
    Signal \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.WriteEnable\: boolean := false;
    Signal \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32).number.parameter.0\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Started.0\: boolean := false;
    Signal \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._Started\: boolean := false;
    Signal \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Finished.0\: boolean := false;
    Signal \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32).return.0\: boolean;
    -- System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 declarations end


    -- System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 declarations start
    -- State machine states:
    type \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._States\ is (
        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_0\, 
        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_1\, 
        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_2\, 
        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_3\, 
        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_4\, 
        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_5\, 
        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_6\, 
        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_7\, 
        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_8\, 
        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_9\, 
        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_10\, 
        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_11\, 
        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_12\);
    -- Signals:
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._Finished\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.CellIndex\: signed(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.DataOut\: std_logic_vector(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.WriteEnable\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.0\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.0\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.1\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.1\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.2\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.2\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.3\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.3\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.4\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.4\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.5\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.5\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.6\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.6\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.7\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.7\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.8\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.8\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.9\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.9\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.10\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.10\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.11\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.11\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.12\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.12\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.13\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.13\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.14\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.14\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.15\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.15\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.16\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.16\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.17\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.17\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.18\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.18\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.19\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.19\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.20\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.20\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.21\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.21\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.22\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.22\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.23\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.23\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.24\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.24\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.25\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.25\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.26\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.26\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.27\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.27\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.28\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.28\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.29\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.29\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.30\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.30\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.31\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.31\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.32\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.32\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.33\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.33\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.34\: unsigned(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.34\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._Started\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.0\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.1\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.2\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.3\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.4\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.5\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.6\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.7\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.8\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.9\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.10\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.11\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.12\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.13\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.14\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.15\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.16\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.17\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.18\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.19\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.20\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.21\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.22\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.23\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.24\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.25\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.26\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.27\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.28\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.29\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.30\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.31\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.32\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.33\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.34\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.0\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.1\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.2\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.3\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.4\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.5\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.6\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.7\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.8\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.9\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.10\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.11\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.12\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.13\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.14\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.15\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.16\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.17\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.18\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.19\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.20\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.21\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.22\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.23\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.24\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.25\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.26\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.27\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.28\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.29\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.30\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.31\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.32\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.33\: boolean;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.34\: boolean;
    -- System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberInternal(System.UInt32).0 declarations start
    -- State machine states:
    type \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._States\ is (
        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_0\, 
        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_1\, 
        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_2\, 
        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_3\, 
        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_4\, 
        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_5\, 
        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_6\, 
        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_7\, 
        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_8\);
    -- Signals:
    Signal \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Finished\: boolean := false;
    Signal \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.return\: boolean;
    Signal \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Started\: boolean := false;
    Signal \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.number.parameter\: unsigned(31 downto 0);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberInternal(System.UInt32).0 declarations end


    -- System.Void Hast::ExternalInvocationProxy() declarations start
    -- Signals:
    Signal \FinishedInternal\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory)._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumberAsync(SimpleMemory)._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().PrimeCalculator::ArePrimeNumbers(SimpleMemory)._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory)._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory)._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumberAsync(SimpleMemory)._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().PrimeCalculator::ArePrimeNumbers(SimpleMemory)._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory)._Finished.0\: boolean := false;
    -- System.Void Hast::ExternalInvocationProxy() declarations end


    -- \System.Void Hast::InternalInvocationProxy()._RunningStates\ declarations start
    type \Hast::InternalInvocationProxy()._RunningStates\ is (
        WaitingForStarted, 
        WaitingForFinished, 
        AfterFinished);
    -- \System.Void Hast::InternalInvocationProxy()._RunningStates\ declarations end

begin 

    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).0 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).0 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).1 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).1 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).2 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).2 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).3 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).3 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).4 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).4 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).5 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).5 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).6 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).6 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).7 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).7 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).8 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).8 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).9 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).9 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).10 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).10 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).11 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).11 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).12 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).12 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).13 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).13 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).14 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).14 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).15 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).15 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).16 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).16 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).17 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).17 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).18 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).18 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).19 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).19 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).20 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).20 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).21 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).21 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).22 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).22 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).23 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).23 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).24 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).24 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).25 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).25 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).26 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).26 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).27 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).27 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).28 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).28 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).29 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).29 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).30 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).30 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).31 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).31 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).32 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).32 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).33 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).33 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).34 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.numberObject\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.flag\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.result\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.numberObject.parameter\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.num3\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object).34 state machine end


    -- System.Void Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumber(Hast.Transformer.SimpleMemory.SimpleMemory).0 state machine start
    \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State\: \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._States\ := \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_0\;
        Variable \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.number\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Finished\ <= false;
                \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.WriteEnable\ <= false;
                \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Started.0\ <= false;
                \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State\ := \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_0\;
            else 
                case \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State\ is 
                    when \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Started\ = true) then 
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State\ := \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Started\ = true) then 
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Finished\ <= true;
                        else 
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Finished\ <= false;
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State\ := \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_2\ => 
                        -- Begin SimpleMemory read.
                        \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.CellIndex\ <= resize(to_signed(0, 32), 32);
                        \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.ReadEnable\ <= true;
                        \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State\ := \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_3\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.number\ := ConvertStdLogicVectorToUInt32(\DataIn\);
                            -- Starting state machine invocation for the following method: System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberInternal(System.UInt32)
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32).number.parameter.0\ <= \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.number\;
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Started.0\ <= true;
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State\ := \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_4\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberInternal(System.UInt32)
                        if (\PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Started.0\ = \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Finished.0\) then 
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Started.0\ <= false;
                            -- Begin SimpleMemory write.
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.CellIndex\ <= resize(to_signed(0, 32), 32);
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.WriteEnable\ <= true;
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.DataOut\ <= ConvertBooleanToStdLogicVector(\PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32).return.0\);
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State\ := \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_5\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\WritesDone\ = true) then 
                            -- SimpleMemory write finished.
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.WriteEnable\ <= false;
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State\ := \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumber(Hast.Transformer.SimpleMemory.SimpleMemory).0 state machine end


    -- System.Threading.Tasks.Task Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberAsync(Hast.Transformer.SimpleMemory.SimpleMemory).0 state machine start
    \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State\: \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._States\ := \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State_0\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._Finished\ <= false;
                \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.PrimeCalculator::IsPrimeNumber(SimpleMemory)._Started.0\ <= false;
                \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State\ := \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State_0\;
            else 
                case \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State\ is 
                    when \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._Started\ = true) then 
                            \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State\ := \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._Started\ = true) then 
                            \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._Finished\ <= true;
                        else 
                            \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._Finished\ <= false;
                            \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State\ := \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State_2\ => 
                        -- Starting state machine invocation for the following method: System.Void Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumber(Hast.Transformer.SimpleMemory.SimpleMemory)
                        \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.PrimeCalculator::IsPrimeNumber(SimpleMemory)._Started.0\ <= true;
                        \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State\ := \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumber(Hast.Transformer.SimpleMemory.SimpleMemory)
                        if (\PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.PrimeCalculator::IsPrimeNumber(SimpleMemory)._Started.0\ = \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.PrimeCalculator::IsPrimeNumber(SimpleMemory)._Finished.0\) then 
                            \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.PrimeCalculator::IsPrimeNumber(SimpleMemory)._Started.0\ <= false;
                            \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State\ := \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Threading.Tasks.Task Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberAsync(Hast.Transformer.SimpleMemory.SimpleMemory).0 state machine end


    -- System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 state machine start
    \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State\: \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._States\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_0\;
        Variable \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.num2\: signed(31 downto 0);
        Variable \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.number\: unsigned(31 downto 0);
        Variable \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.0\: boolean;
        Variable \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.2\: signed(31 downto 0);
        Variable \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.3\: signed(31 downto 0);
        Variable \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.4\: signed(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._Finished\ <= false;
                \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.WriteEnable\ <= false;
                \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Started.0\ <= false;
                \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_0\;
            else 
                case \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State\ is 
                    when \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._Started\ = true) then 
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._Started\ = true) then 
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._Finished\ <= true;
                        else 
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._Finished\ <= false;
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_2\ => 
                        -- Begin SimpleMemory read.
                        \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.CellIndex\ <= resize(to_signed(0, 32), 32);
                        \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\ <= true;
                        \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_3\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.num\ := ConvertStdLogicVectorToUInt32(\DataIn\);
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.num2\ := to_signed(0, 32);
                            -- Starting a while loop.
                            -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.0\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.num2\ < signed((\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.num\));
                            if (\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.0\) then 
                                \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_4\;
                            else 
                                \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_5\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_4\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_3\.
                        -- The while loop's condition:
                        \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.1\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.num2\ < signed((\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.num\));
                        if (\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.1\) then 
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.2\ := to_signed(1, 32) + \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.num2\;
                            -- Begin SimpleMemory read.
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.CellIndex\ <= resize(\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.2\, 32);
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\ <= true;
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_6\;
                        else 
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_5\ => 
                        -- State after the while loop which was started in state \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_3\.
                        \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_6\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.number\ := ConvertStdLogicVectorToUInt32(\DataIn\);
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.3\ := to_signed(1, 32) + \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.num2\;
                            -- Starting state machine invocation for the following method: System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberInternal(System.UInt32)
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32).number.parameter.0\ <= \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.number\;
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Started.0\ <= true;
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_7\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberInternal(System.UInt32)
                        if (\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Started.0\ = \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Finished.0\) then 
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Started.0\ <= false;
                            -- Begin SimpleMemory write.
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.CellIndex\ <= resize(\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.3\, 32);
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.WriteEnable\ <= true;
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.DataOut\ <= ConvertBooleanToStdLogicVector(\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32).return.0\);
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_8\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_8\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\WritesDone\ = true) then 
                            -- SimpleMemory write finished.
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.WriteEnable\ <= false;
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.4\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.num2\ + to_signed(1, 32);
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.num2\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.4\;
                            -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_3\ if the loop wasn't exited with a state change.
                            if (\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State\ = \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_8\) then 
                                \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_4\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 state machine end


    -- System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 state machine start
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\: \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._States\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_0\;
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\: boolean_Array(0 to 34);
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num2\: signed(31 downto 0);
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.i\: signed(31 downto 0);
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\: unsigned(31 downto 0);
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.arg_5D_1\: signed(31 downto 0);
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.j\: signed(31 downto 0);
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.0\: boolean;
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.3\: boolean;
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.4\: signed(31 downto 0);
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.5\: signed(31 downto 0);
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).invocationIndex\: integer range 0 to 34 := 0;
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.6\: signed(31 downto 0);
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.7\: boolean;
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.8\: boolean;
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.9\: signed(31 downto 0);
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.10\: signed(31 downto 0);
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.11\: signed(31 downto 0);
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.12\: signed(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._Finished\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.WriteEnable\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.0\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.1\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.2\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.3\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.4\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.5\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.6\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.7\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.8\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.9\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.10\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.11\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.12\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.13\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.14\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.15\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.16\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.17\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.18\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.19\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.20\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.21\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.22\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.23\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.24\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.25\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.26\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.27\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.28\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.29\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.30\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.31\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.32\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.33\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.34\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_0\;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).invocationIndex\ := 0;
            else 
                case \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ is 
                    when \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._Started\ = true) then 
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._Started\ = true) then 
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._Finished\ <= true;
                        else 
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._Finished\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_2\ => 
                        -- Begin SimpleMemory read.
                        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.CellIndex\ <= resize(to_signed(0, 32), 32);
                        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\ <= true;
                        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_3\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num\ := ConvertStdLogicVectorToUInt32(\DataIn\);
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\ := (others => false);
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num2\ := to_signed(0, 32);
                            -- Starting a while loop.
                            -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.0\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num2\ < signed((\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num\));
                            if (\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.0\) then 
                                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_4\;
                            else 
                                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_5\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_4\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_3\.
                        -- The while loop's condition:
                        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.1\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num2\ < signed((\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num\));
                        if (\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.1\) then 
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.i\ := to_signed(0, 32);
                            -- Starting a while loop.
                            -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.2\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.i\ < to_signed(35, 32);
                            if (\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.2\) then 
                                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_6\;
                            else 
                                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_7\;
                            end if;
                        else 
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_5\ => 
                        -- State after the while loop which was started in state \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_3\.
                        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_6\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_4\.
                        -- The while loop's condition:
                        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.3\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.i\ < to_signed(35, 32);
                        if (\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.3\) then 
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.4\ := to_signed(1, 32) + \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num2\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.5\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.4\ + \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.i\;
                            -- Begin SimpleMemory read.
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.CellIndex\ <= resize(\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.5\, 32);
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\ <= true;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_8\;
                        else 
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,3
                    when \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_7\ => 
                        -- State after the while loop which was started in state \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_4\.
                        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_9\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_8\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\ := ConvertStdLogicVectorToUInt32(\DataIn\);
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.arg_5D_1\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.i\;
                            -- Starting state machine invocation for the following method: System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object)
                            case \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).invocationIndex\ is 
                                when 0 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.0\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.0\ <= true;
                                when 1 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.1\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.1\ <= true;
                                when 2 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.2\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.2\ <= true;
                                when 3 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.3\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.3\ <= true;
                                when 4 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.4\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.4\ <= true;
                                when 5 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.5\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.5\ <= true;
                                when 6 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.6\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.6\ <= true;
                                when 7 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.7\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.7\ <= true;
                                when 8 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.8\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.8\ <= true;
                                when 9 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.9\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.9\ <= true;
                                when 10 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.10\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.10\ <= true;
                                when 11 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.11\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.11\ <= true;
                                when 12 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.12\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.12\ <= true;
                                when 13 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.13\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.13\ <= true;
                                when 14 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.14\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.14\ <= true;
                                when 15 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.15\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.15\ <= true;
                                when 16 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.16\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.16\ <= true;
                                when 17 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.17\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.17\ <= true;
                                when 18 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.18\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.18\ <= true;
                                when 19 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.19\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.19\ <= true;
                                when 20 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.20\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.20\ <= true;
                                when 21 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.21\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.21\ <= true;
                                when 22 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.22\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.22\ <= true;
                                when 23 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.23\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.23\ <= true;
                                when 24 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.24\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.24\ <= true;
                                when 25 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.25\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.25\ <= true;
                                when 26 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.26\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.26\ <= true;
                                when 27 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.27\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.27\ <= true;
                                when 28 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.28\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.28\ <= true;
                                when 29 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.29\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.29\ <= true;
                                when 30 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.30\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.30\ <= true;
                                when 31 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.31\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.31\ <= true;
                                when 32 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.32\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.32\ <= true;
                                when 33 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.33\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.33\ <= true;
                                when 34 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.34\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.34\ <= true;
                            end case;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).invocationIndex\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).invocationIndex\ + 1;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.6\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.i\ + to_signed(1, 32);
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.i\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.6\;
                            -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_4\ if the loop wasn't exited with a state change.
                            if (\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_8\) then 
                                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_6\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_9\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object)
                        if (\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.1\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.1\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.2\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.2\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.3\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.3\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.4\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.4\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.5\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.5\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.6\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.6\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.7\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.7\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.8\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.8\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.9\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.9\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.10\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.10\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.11\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.11\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.12\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.12\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.13\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.13\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.14\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.14\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.15\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.15\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.16\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.16\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.17\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.17\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.18\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.18\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.19\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.19\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.20\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.20\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.21\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.21\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.22\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.22\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.23\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.23\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.24\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.24\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.25\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.25\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.26\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.26\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.27\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.27\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.28\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.28\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.29\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.29\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.30\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.30\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.31\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.31\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.32\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.32\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.33\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.33\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.34\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.34\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.0\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.0\) then 
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.0\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.1\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.2\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.3\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.4\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.5\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.6\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.7\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.8\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.9\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.10\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.11\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.12\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.13\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.14\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.15\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.16\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.17\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.18\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.19\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.20\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.21\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.22\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.23\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.24\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.25\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.26\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.27\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.28\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.29\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.30\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.31\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.32\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.33\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.34\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).invocationIndex\ := 0;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(0) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.0\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(1) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.1\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(2) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.2\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(3) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.3\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(4) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.4\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(5) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.5\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(6) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.6\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(7) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.7\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(8) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.8\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(9) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.9\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(10) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.10\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(11) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.11\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(12) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.12\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(13) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.13\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(14) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.14\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(15) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.15\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(16) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.16\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(17) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.17\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(18) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.18\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(19) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.19\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(20) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.20\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(21) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.21\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(22) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.22\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(23) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.23\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(24) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.24\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(25) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.25\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(26) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.26\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(27) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.27\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(28) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.28\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(29) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.29\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(30) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.30\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(31) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.31\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(32) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.32\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(33) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.33\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(34) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.34\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.j\ := to_signed(0, 32);
                            -- Starting a while loop.
                            -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.7\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.j\ < to_signed(35, 32);
                            if (\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.7\) then 
                                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_10\;
                            else 
                                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_11\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_10\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_9\.
                        -- The while loop's condition:
                        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.8\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.j\ < to_signed(35, 32);
                        if (\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.8\) then 
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.9\ := to_signed(1, 32) + \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num2\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.10\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.9\ + \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.j\;
                            -- Begin SimpleMemory write.
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.CellIndex\ <= resize(\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.10\, 32);
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.WriteEnable\ <= true;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.DataOut\ <= ConvertBooleanToStdLogicVector(\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(to_integer(\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.j\)));
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_12\;
                        else 
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_11\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,3
                    when \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_11\ => 
                        -- State after the while loop which was started in state \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_9\.
                        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.12\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num2\ + to_signed(35, 32);
                        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num2\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.12\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_3\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_11\) then 
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_12\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\WritesDone\ = true) then 
                            -- SimpleMemory write finished.
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.WriteEnable\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.11\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.j\ + to_signed(1, 32);
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.j\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.11\;
                            -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_9\ if the loop wasn't exited with a state change.
                            if (\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_12\) then 
                                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_10\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberInternal(System.UInt32).0 state machine start
    \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\: \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._States\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_0\;
        Variable \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.number\: unsigned(31 downto 0);
        Variable \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.num\: unsigned(31 downto 0);
        Variable \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.num2\: unsigned(31 downto 0);
        Variable \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.flag\: boolean;
        Variable \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.result\: boolean;
        Variable \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.0\: unsigned(31 downto 0);
        Variable \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.1\: boolean;
        Variable \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.2\: boolean;
        Variable \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.3\: unsigned(31 downto 0);
        Variable \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.4\: boolean;
        Variable \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.5\: unsigned(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Finished\ <= false;
                \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_0\;
                \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ is 
                    when \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Started\ = true) then 
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Started\ = true) then 
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Finished\ <= true;
                        else 
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Finished\ <= false;
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_2\ => 
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.number\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.number.parameter\;
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.0\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.number\ / to_unsigned(2, 32);
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.num\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.0\;
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.num2\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.1\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.num2\ <= \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.num\;
                        if (\PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.1\) then 
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_3\;
                        else 
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,2
                    when \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.2\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.num2\ <= \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.num\;
                        if (\PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.2\) then 
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_5\;
                        else 
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_2\.
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.result\ := True;
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.return\ <= \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.result\;
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.3\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.number\ mod \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.num2\;
                        if (\PrimeCalculator::IsPrimeNumberInternal(UInt32).0.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_6\;
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_6\ => 
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.4\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.flag\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_8\ and ends in state \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_7\.

                        if (\PrimeCalculator::IsPrimeNumberInternal(UInt32).0.flag\) then 
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_6\.
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.5\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.num2\ + to_unsigned(1, 32);
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.num2\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ = \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_7\) then 
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0,1
                    when \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_6\.
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.result\ := False;
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.return\ <= \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.result\;
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_6\.
                        if (\PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ = \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_8\) then 
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberInternal(System.UInt32).0 state machine end


    -- System.Void Hast::ExternalInvocationProxy() start
    \Finished\ <= \FinishedInternal\;
    \Hast::ExternalInvocationProxy()\: process (\Clock\) 
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \FinishedInternal\ <= false;
                \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory)._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumberAsync(SimpleMemory)._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().PrimeCalculator::ArePrimeNumbers(SimpleMemory)._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory)._Started.0\ <= false;
            else 
                if (\Started\ = true and \FinishedInternal\ = false) then 
                    -- Starting the state machine corresponding to the given member ID.
                    case \MemberId\ is 
                        when 0 => 
                            if (\Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory)._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory)._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory)._Started.0\ = \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory)._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory)._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 1 => 
                            if (\Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumberAsync(SimpleMemory)._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumberAsync(SimpleMemory)._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumberAsync(SimpleMemory)._Started.0\ = \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumberAsync(SimpleMemory)._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumberAsync(SimpleMemory)._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 2 => 
                            if (\Hast::ExternalInvocationProxy().PrimeCalculator::ArePrimeNumbers(SimpleMemory)._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().PrimeCalculator::ArePrimeNumbers(SimpleMemory)._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().PrimeCalculator::ArePrimeNumbers(SimpleMemory)._Started.0\ = \Hast::ExternalInvocationProxy().PrimeCalculator::ArePrimeNumbers(SimpleMemory)._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().PrimeCalculator::ArePrimeNumbers(SimpleMemory)._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 3 => 
                            if (\Hast::ExternalInvocationProxy().PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory)._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory)._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory)._Started.0\ = \Hast::ExternalInvocationProxy().PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory)._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory)._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when others => 
                            null;
                    end case;
                else 
                    -- Waiting for Started to be pulled back to zero that signals the framework noting the finish.
                    if (\Started\ = false and \FinishedInternal\ = true) then 
                        \FinishedInternal\ <= false;
                    end if;
                end if;
            end if;
        end if;
    end process;
    -- System.Void Hast::ExternalInvocationProxy() end


    -- System.Void Hast::InternalInvocationProxy().System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberInternal(System.UInt32) start
    \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Started\: boolean := false;
        Variable \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumberInternal(UInt32).0.justFinished\: boolean;
        Variable \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumber(SimpleMemory).0.runningIndex.0\: integer range 0 to 0;
        Variable \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumber(SimpleMemory).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.runningIndex.0\: integer range 0 to 0;
        Variable \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Started\ := false;
                \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumber(SimpleMemory).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.runningState.0\ := WaitingForStarted;
                \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Finished.0\ <= false;
                \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Finished.0\ <= false;
            else 

                -- Temporary Started variables are needed in place of the original signals so inside the proxy it's immediately visible if an instance is already started.
                \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Started\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Started\;


                -- JustFinished states should be only kept for one clock cycle, since they are used not to immediately restart a state machine once it finished.
                \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumberInternal(UInt32).0.justFinished\ := false;


                -- Invocation handler #0 out of 1 corresponding to System.Void Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumber(Hast.Transformer.SimpleMemory.SimpleMemory).0
                case \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumber(SimpleMemory).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Started.0\) then 
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Finished.0\ <= false;
                            if (\Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Started\ = false and \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumberInternal(UInt32).0.justFinished\ = false) then 
                                \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumber(SimpleMemory).0.runningState.0\ := WaitingForFinished;
                                \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumber(SimpleMemory).0.runningIndex.0\ := 0;
                                \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Started\ := true;
                                \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.number.parameter\ <= \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32).number.parameter.0\;
                            end if;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumber(SimpleMemory).0.runningIndex.0\ is 
                            when 0 => 
                                if (\PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumber(SimpleMemory).0.runningState.0\ := AfterFinished;
                                    \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Finished.0\ <= true;
                                    \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Started\ := false;
                                    \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumberInternal(UInt32).0.justFinished\ := true;
                                    \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32).return.0\ <= \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumber(SimpleMemory).0.runningState.0\ := WaitingForStarted;
                            case \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumber(SimpleMemory).0.runningIndex.0\ is 
                                when 0 => 
                                    \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Finished.0\ <= false;
                            end case;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0
                case \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Started.0\) then 
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Finished.0\ <= false;
                            if (\Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Started\ = false and \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumberInternal(UInt32).0.justFinished\ = false) then 
                                \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.runningState.0\ := WaitingForFinished;
                                \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.runningIndex.0\ := 0;
                                \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Started\ := true;
                                \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.number.parameter\ <= \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32).number.parameter.0\;
                            end if;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.runningIndex.0\ is 
                            when 0 => 
                                if (\PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.runningState.0\ := AfterFinished;
                                    \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Finished.0\ <= true;
                                    \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Started\ := false;
                                    \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumberInternal(UInt32).0.justFinished\ := true;
                                    \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32).return.0\ <= \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.runningState.0\ := WaitingForStarted;
                            case \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.runningIndex.0\ is 
                                when 0 => 
                                    \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Finished.0\ <= false;
                            end case;
                        end if;
                end case;


                -- Writing Started variable values back to signals.
                \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Started\ <= \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Started\;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberInternal(System.UInt32) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumber(Hast.Transformer.SimpleMemory.SimpleMemory) start
    \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Started\: boolean := false;
        Variable \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumber(SimpleMemory).0.justFinished\: boolean;
        Variable \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.runningIndex.0\: integer range 0 to 0;
        Variable \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).Hast::ExternalInvocationProxy().runningIndex.0\: integer range 0 to 0;
        Variable \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).Hast::ExternalInvocationProxy().runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Started\ := false;
                \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).Hast::ExternalInvocationProxy().runningState.0\ := WaitingForStarted;
                \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.PrimeCalculator::IsPrimeNumber(SimpleMemory)._Finished.0\ <= false;
                \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory)._Finished.0\ <= false;
            else 

                -- Temporary Started variables are needed in place of the original signals so inside the proxy it's immediately visible if an instance is already started.
                \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Started\ := \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Started\;


                -- JustFinished states should be only kept for one clock cycle, since they are used not to immediately restart a state machine once it finished.
                \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumber(SimpleMemory).0.justFinished\ := false;


                -- Invocation handler #0 out of 1 corresponding to System.Threading.Tasks.Task Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberAsync(Hast.Transformer.SimpleMemory.SimpleMemory).0
                case \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.PrimeCalculator::IsPrimeNumber(SimpleMemory)._Started.0\) then 
                            \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.PrimeCalculator::IsPrimeNumber(SimpleMemory)._Finished.0\ <= false;
                            if (\Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Started\ = false and \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumber(SimpleMemory).0.justFinished\ = false) then 
                                \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.runningState.0\ := WaitingForFinished;
                                \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.runningIndex.0\ := 0;
                                \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Started\ := true;
                            end if;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.runningIndex.0\ is 
                            when 0 => 
                                if (\PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.runningState.0\ := AfterFinished;
                                    \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.PrimeCalculator::IsPrimeNumber(SimpleMemory)._Finished.0\ <= true;
                                    \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Started\ := false;
                                    \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumber(SimpleMemory).0.justFinished\ := true;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.PrimeCalculator::IsPrimeNumber(SimpleMemory)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.runningState.0\ := WaitingForStarted;
                            case \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.runningIndex.0\ is 
                                when 0 => 
                                    \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.PrimeCalculator::IsPrimeNumber(SimpleMemory)._Finished.0\ <= false;
                            end case;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Void Hast::ExternalInvocationProxy()
                case \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).Hast::ExternalInvocationProxy().runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory)._Started.0\) then 
                            \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory)._Finished.0\ <= false;
                            if (\Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Started\ = false and \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumber(SimpleMemory).0.justFinished\ = false) then 
                                \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).Hast::ExternalInvocationProxy().runningState.0\ := WaitingForFinished;
                                \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).Hast::ExternalInvocationProxy().runningIndex.0\ := 0;
                                \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Started\ := true;
                            end if;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).Hast::ExternalInvocationProxy().runningIndex.0\ is 
                            when 0 => 
                                if (\PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).Hast::ExternalInvocationProxy().runningState.0\ := AfterFinished;
                                    \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory)._Finished.0\ <= true;
                                    \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Started\ := false;
                                    \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumber(SimpleMemory).0.justFinished\ := true;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).Hast::ExternalInvocationProxy().runningState.0\ := WaitingForStarted;
                            case \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).Hast::ExternalInvocationProxy().runningIndex.0\ is 
                                when 0 => 
                                    \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory)._Finished.0\ <= false;
                            end case;
                        end if;
                end case;


                -- Writing Started variable values back to signals.
                \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Started\ <= \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Started\;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumber(Hast.Transformer.SimpleMemory.SimpleMemory) end


    -- System.Void Hast::InternalInvocationProxy().System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object) start
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#0):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.0\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.0\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.0\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.0\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).0.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#1):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.1\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.1\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.1\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.1\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).1.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#2):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.2\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.2\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.2\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.2\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).2.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#3):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.3\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.3\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).3.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#4):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.4\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.4\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.4\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.4\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).4.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#5):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.5\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.5\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.5\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.5\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).5.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#6):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.6\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.6\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.6\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.6\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).6.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#7):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.7\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.7\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.7\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.7\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).7.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#8):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.8\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.8\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.8\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.8\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).8.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#9):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.9\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.9\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.9\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.9\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).9.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#10):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.10\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.10\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.10\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.10\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).10.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#11):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.11\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.11\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.11\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.11\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).11.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#12):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.12\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.12\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.12\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.12\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).12.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#13):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.13\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.13\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.13\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.13\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).13.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#14):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.14\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.14\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.14\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.14\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).14.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#15):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.15\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.15\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.15\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.15\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).15.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#16):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.16\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.16\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.16\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.16\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).16.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#17):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.17\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.17\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.17\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.17\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).17.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#18):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.18\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.18\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.18\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.18\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).18.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#19):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.19\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.19\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.19\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.19\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).19.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#20):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.20\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.20\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.20\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.20\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).20.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#21):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.21\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.21\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.21\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.21\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).21.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#22):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.22\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.22\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.22\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.22\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).22.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#23):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.23\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.23\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.23\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.23\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).23.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#24):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.24\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.24\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.24\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.24\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).24.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#25):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.25\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.25\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.25\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.25\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).25.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#26):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.26\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.26\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.26\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.26\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).26.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#27):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.27\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.27\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.27\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.27\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).27.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#28):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.28\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.28\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.28\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.28\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).28.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#29):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.29\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.29\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.29\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.29\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).29.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#30):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.30\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.30\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.30\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.30\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).30.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#31):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.31\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.31\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.31\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.31\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).31.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#32):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.32\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.32\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.32\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.32\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).32.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#33):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.33\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.33\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.33\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.33\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).33.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory).0 (#34):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Started.34\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.numberObject.parameter\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).numberObject.parameter.34\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object)._Finished.34\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).return.34\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(Object).34.return\;
    -- System.Void Hast::InternalInvocationProxy().System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.Object) end


    -- System.Void Hast::InternalInvocationProxy().System.Threading.Tasks.Task Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberAsync(Hast.Transformer.SimpleMemory.SimpleMemory) start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._Started\ <= \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumberAsync(SimpleMemory)._Started.0\;
    \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumberAsync(SimpleMemory)._Finished.0\ <= \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Threading.Tasks.Task Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberAsync(Hast.Transformer.SimpleMemory.SimpleMemory) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory) start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._Started\ <= \Hast::ExternalInvocationProxy().PrimeCalculator::ArePrimeNumbers(SimpleMemory)._Started.0\;
    \Hast::ExternalInvocationProxy().PrimeCalculator::ArePrimeNumbers(SimpleMemory)._Finished.0\ <= \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory) start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._Started\ <= \Hast::ExternalInvocationProxy().PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory)._Started.0\;
    \Hast::ExternalInvocationProxy().PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory)._Finished.0\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.SimpleMemory.SimpleMemory) end


    -- System.Void Hast::SimpleMemoryOperationProxy() start
    \CellIndex\ <= to_integer(\PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.CellIndex\) when \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.ReadEnable\ or \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.WriteEnable\ else to_integer(\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.CellIndex\) when \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\ or \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.WriteEnable\ else to_integer(\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.CellIndex\) when \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\ or \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.WriteEnable\ else 0;
    \DataOut\ <= \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.DataOut\ when \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.WriteEnable\ else \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.DataOut\ when \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.WriteEnable\ else \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.DataOut\ when \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.WriteEnable\ else "00000000000000000000000000000000";
    \ReadEnable\ <= \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\ or \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\ or \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.ReadEnable\;
    \WriteEnable\ <= \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.WriteEnable\ or \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.WriteEnable\ or \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.WriteEnable\;
    -- System.Void Hast::SimpleMemoryOperationProxy() end

end Imp;
